library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.PhoenixPackage.all;

package TablePackage is

constant NREG : integer := 6;
constant MEMORY_SIZE : integer := NREG;

type memory is array (0 to MEMORY_SIZE-1) of reg26;
type tables is array (0 to NROT-1) of memory;

constant TAB: tables :=(
 -- Router 00
(("10000000000010000010000100"),
("10000000100000100010000001"),
("00000000000000000000000000"),
("00000000000000000000000000"),
("00000000000000000000000000"),
("00000000000000000000000000")
),
 -- Router 01
(("11100000100000100000100001"),
("11001000000100100010000100"),
("10101000000000000000001000"),
("00000000000000000000000000"),
("00000000000000000000000000"),
("00000000000000000000000000")
),
 -- Router 02
(("10101000000000000000101000"),
("11001000000110100010000100"),
("11100000100000100001000001"),
("00000000000000000000000000"),
("00000000000000000000000000"),
("00000000000000000000000000")
),
 -- Router 03
(("11100000100110010001100001"),
("11001000001000010010000100"),
("11100001100110100010000001"),
("10101000000000100001001000"),
("00000000000000000000000000"),
("00000000000000000000000000")
),
 -- Router 04
(("11000000101000010010000001"),
("10000001100000100010001001"),
("10001000000000010001101000"),
("00000000000000000000000000"),
("00000000000000000000000000"),
("00000000000000000000000000")
),
 -- Router 10
(("10101000000000000000000010"),
("10010000000010001010000100"),
("10010001000000100010000001"),
("00000000000000000000000000"),
("00000000000000000000000000"),
("00000000000000000000000000")
),
 -- Router 11
(("10111000000000001000001000"),
("11001000000000000000100010"),
("11110001000000100000100001"),
("11001000000100100010000100"),
("00000000000000000000000000"),
("00000000000000000000000000")
),
 -- Router 12
(("11110001000100010001000001"),
("10111000000000000000001000"),
("11001000000000000010000010"),
("11110001100100100010000001"),
("11001000100110100010000100"),
("10111000100000100000101000")
),
 -- Router 13
(("11110001000110010001100001"),
("11011000101000010010000100"),
("11110001100110100010000001"),
("11101000000000000010000010"),
("10111000100000100001001000"),
("00000000000000000000000000")
),
 -- Router 14
(("10001000001000000010000010"),
("10000001100000100010001001"),
("10001000000000010001101000"),
("11010001000000100010000001"),
("00000000000000000000000000"),
("00000000000000000000000000")
),
 -- Router 20
(("10101000000000001000000010"),
("10010001100000100010000001"),
("10010000000010010010000100"),
("00000000000000000000000000"),
("00000000000000000000000000"),
("00000000000000000000000000")
),
 -- Router 21
(("10111000000000010000001000"),
("11110001100000100000100001"),
("11001000000000001000100010"),
("11001000000100100010000100"),
("00000000000000000000000000"),
("00000000000000000000000000")
),
 -- Router 22
(("10111001000000010000101000"),
("10111000000000001000001000"),
("11001000000000001001000010"),
("11110001100000100010000001"),
("11001000000110100010000100"),
("00000000000000000000000000")
),
 -- Router 23
(("10111000000000001000001000"),
("11001000001000010010000100"),
("11110001100110100010000001"),
("11001000000000001001100010"),
("10111001000000100001001000"),
("00000000000000000000000000")
),
 -- Router 24
(("10010001000000010001101000"),
("10010001100000100010001000"),
("11000000000000001010000010"),
("00000000000000000000000000"),
("00000000000000000000000000"),
("00000000000000000000000000")
),
 -- Router 30
(("10101000000000010000000010"),
("10010010000000100010000001"),
("10010000000010011010000100"),
("00000000000000000000000000"),
("00000000000000000000000000"),
("00000000000000000000000000")
),
 -- Router 31
(("11110010000000100000100001"),
("10111000000000011000001000"),
("11001000000000010000100010"),
("11001000000100100010000100"),
("00000000000000000000000000"),
("00000000000000000000000000")
),
 -- Router 32
(("11011001100110011010000100"),
("11110010000100100010000001"),
("10111001100000100000101000"),
("11101000000000010010000010"),
("00000000000000000000000000"),
("00000000000000000000000000")
),
 -- Router 33
(("11011001101000011010000100"),
("11110010000110100010000001"),
("10101000000110010010000010"),
("10101000000000100001001000"),
("00000000000000000000000000"),
("00000000000000000000000000")
),
 -- Router 34
(("10000001100000011001101000"),
("10000010000000100010000001"),
("10000000000000010010001000"),
("00000000000000000000000000"),
("00000000000000000000000000"),
("00000000000000000000000000")
),
 -- Router 40
(("10010000000010100010000100"),
("10100000000000011000000010"),
("00000000000000000000000000"),
("00000000000000000000000000"),
("00000000000000000000000000"),
("00000000000000000000000000")
),
 -- Router 41
(("10110000000000100000001000"),
("11000000000000011000100010"),
("11000000000100100010000100"),
("00000000000000000000000000"),
("00000000000000000000000000"),
("00000000000000000000000000")
),
 -- Router 42
(("11010010000110100010000100"),
("10110010000000100000101000"),
("11100000000000011010000010"),
("00000000000000000000000000"),
("00000000000000000000000000"),
("00000000000000000000000000")
),
 -- Router 43
(("11010001101000100010000100"),
("10100000000110011010000010"),
("10100000000000100001001000"),
("00000000000000000000000000"),
("00000000000000000000000000"),
("00000000000000000000000000")
),
 -- Router 44
(("11000001101000011010000010"),
("10010000000000010010001000"),
("10010001100000100001101000"),
("00000000000000000000000000"),
("00000000000000000000000000"),
("00000000000000000000000000")
)
);
end TablePackage;

package body TablePackage is
end TablePackage;
